package Types is  

type ULA_OP is (AND_OP, OR_OP, ADD_OP, ADDU_OP,
                SUB_OP, SUBU_OP, SLT_OP, SLTU_OP, 
                NOR_OP, XOR_OP, SLL_OP, SRL_OP,  
                SRA_OP, RTR_OP, RTL_OP); 
end Types;
